library IEEE; use IEEE.std_logic_1164.all;

entity f_system is

  port ( x1, x2, x3, x4: in std_logic;

         y1, y2, y3, y4: out std_logic );

end entity f_system;
